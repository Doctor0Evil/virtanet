module noc_interconnect (/* inputs, outputs */);
  // Reconfigurable interconnect fabric for spike routing
endmodule
