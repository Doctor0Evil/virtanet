module ccm_control_unit (/* inputs, outputs */);
  // AXI-Lite slave interface, interrupt controller, PMU, DMA controller logic
endmodule
