module npu_core (/* inputs, outputs */);
  // Leaky Integrate-and-Fire neuron model, STDP logic
endmodule
