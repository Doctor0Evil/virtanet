module on_chip_memory (/* inputs, outputs */);
  // High-speed SRAM for weights, NPU states, spike buffers
endmodule
