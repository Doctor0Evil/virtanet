module top_ccm (/* inputs, outputs */);
  // Instantiation of CCU, NPU Array, NoC, OCM
endmodule
